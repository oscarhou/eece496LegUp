library ieee;
use ieee.std_logic_1164.all;
library work;
use work.sha3_types.all;

ENTITY theta IS
	PORT(inData: in row);
END theta;