-- Chi step
library ieee;
use ieee.std_logic_1164.all;

ENTITY chi IS
end chi;