--Iota step
library ieee;	
use ieee.std_logic_1164.all;