library ieee;
use ieee.std_logic_1164.all;
library work;
use work.sha3_types.all;

ENTITY sha3 IS
PORT(inputState :in lane);
END sha3;

ARCHITECTURE shaArch OF sha3 IS
BEGIN
END shaArch;