-- Rho and Pi steps of the round function
library ieee;
use ieee.std_logic_1164.all;